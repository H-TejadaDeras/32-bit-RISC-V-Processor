/* 
 *  Processor Registers
 *
 *  Declares Conventional RISC-V RV32I Registers
 *  Conventional Registers:
 *  x0 - Zero
 *  x1 - ra
 *  ...
 */