/*
 *  RISC-V Processor with RV32I Instructions
 */