/*
 *  Arithmetic Logic Unit
 *  
 *  Computes Addition and Subtraction Operations
 *  Supported Operations:
 *  ...
 */

 