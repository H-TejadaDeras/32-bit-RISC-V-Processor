/*
 *  Instruction Decoder Module
 *  
 *  Decodes RISC-V RV32I Instructions
 *  Implemented Instructions:
 *  ...
 */