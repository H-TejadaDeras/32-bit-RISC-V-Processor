/*
 *  RISC-V Processor with RV32I Instructions
 */

`include "memory.sv"
`include "pc.sv"
`include "registers.sv"
`include "decoder.sv"

module top (
    input logic clk, 
    output logic LED, 
    output logic RGB_R, 
    output logic RGB_G, 
    output logic RGB_B
);
   // variables for controlling LED
    localparam [3:0] INIT       = 4'd0;
    localparam [3:0] RED        = 4'd1;
    localparam [3:0] YELLOW     = 4'd2;
    localparam [3:0] GREEN      = 4'd3;
    localparam [3:0] CYAN       = 4'd4;
    localparam [3:0] BLUE       = 4'd5;
    localparam [3:0] MAGENTA    = 4'd6;
    localparam [21:0] STATE_DWELL_CYCLES = 22'd3000000;


    // values for storing/retriving memory
    logic [2:0] funct3 = 3'b010;
    logic dmem_wren = 1'b0;
    logic [31:0] dmem_address = 31'd0;
    logic [31:0] dmem_data_in = 31'd0;
    logic [31:0] dmem_data_out;
    logic [31:0] imem_address = 31'h1000;
    logic [31:0] imem_data_out;
    logic reset;

    // values for program counter
    logic [1:0] instruction_completed = 1'b1;
    logic [31:0] increment = 32'd4;
    logic [31:0] instruction_output;

    // Variables for reading from a register and writing to register
    logic [31:0] reg_address = 32'h00000002; // Stack Pointer
    logic [31:0] reg_input = 32'h01010101;
    logic        reg_operation = 1'b1;
    logic [31:0] reg_output;
    logic [31:0] tmp;

    // variables for signals
    logic led;
    logic red;
    logic green;
    logic blue;

    // variables for decoder
    logic [6:0]  opcode;
    logic [4:0]  rd;
    logic [2:0]  funct3_out;
    logic [4:0]  rs1;
    logic [4:0]  rs2;
    logic [6:0]  funct7;
    logic [31:0] imm_i;
    logic [31:0] imm_s;
    logic [31:0] imm_b;
    logic [31:0] imm_u;
    logic [31:0] imm_j;
    logic [4:0] index;

    logic [3:0] state = INIT;
    logic [21:0] count = 22'd0;


    program_counter u1 (
        .clk                       (clk), 
        .instruction_completed     (instruction_completed[1:0]),
        .imem_address              (imem_address[31:0]),
        .increment                 (increment[31:0]),
        .instruction               (instruction_output[31:0])
    );

    decoder u2 (
        .clk                       (clk),
        .instruction               (imem_data_out),
        .opcode                    (opcode),
        .rd                        (rd),
        .funct3                    (funct3_out),
        .rs1                       (rs1),
        .rs2                       (rs2),
        .funct7                    (funct7),
        .imm_i                     (imm_i),
        .imm_s                     (imm_s),
        .imm_b                     (imm_b),
        .imm_u                     (imm_u),
        .imm_j                     (imm_j),
        .index                     (index)
    );

    // registers u3 (
    //     .clk                        (clk),
    //     .reg_address                (reg_address[31:0]),
    //     .reg_input                  (reg_input[31:0]),
    //     .reg_operation              (reg_operation),
    //     .reg_output                 (reg_output[31:0])
    // );

    // Testing Code for Register Functions
    // always_ff @(posedge clk) begin
    //     reg_input <= ~reg_input;
    //     // reg_operation <= ~reg_operation;
    // end

    // brad's code for controlling LEDs we can delete it but its here for reference.
    always_ff @(negedge clk) begin
        imem_address <= instruction_output;
        case (state)
            INIT: begin
                dmem_address <= 32'hFFFFFFFC;
                dmem_data_in <= 32'hFFFF0000;
                dmem_wren <= 1'b1;
                count <= STATE_DWELL_CYCLES;
                state <= RED;
            end
            RED: begin
                if (count > 22'd0) begin
                    count <= count - 1;
                end
                else begin
                    dmem_data_in <= 32'hFFFFFF00;
                    count <= STATE_DWELL_CYCLES;
                    state <= YELLOW;
                end
            end
            YELLOW: begin
                if (count > 22'd0) begin
                    count <= count - 1;
                end
                else begin
                    dmem_data_in <= 32'hFF00FF00;
                    count <= STATE_DWELL_CYCLES;
                    state <= GREEN;
                end
            end
            GREEN: begin
                if (count > 22'd0) begin
                    count <= count - 1;
                end
                else begin
                    dmem_data_in <= 32'h0000FFFF;
                    count <= STATE_DWELL_CYCLES;
                    state <= CYAN;
                end
            end
            CYAN: begin
                if (count > 22'd0) begin
                    count <= count - 1;
                end
                else begin
                    dmem_data_in <= 32'h000000FF;
                    count <= STATE_DWELL_CYCLES;
                    state <= BLUE;
                end
            end
            BLUE: begin
                if (count > 22'd0) begin
                    count <= count - 1;
                end
                else begin
                    dmem_data_in <= 32'h00FF00FF;
                    count <= STATE_DWELL_CYCLES;
                    state <= MAGENTA;
                end
            end
            MAGENTA: begin
                if (count > 22'd0) begin
                    count <= count - 1;
                end
                else begin
                    dmem_data_in <= 32'hFFFF0000;
                    count <= STATE_DWELL_CYCLES;
                    state <= RED;
                end
            end
        endcase
    end

    memory #(
        .IMEM_INIT_FILE_PREFIX  ("example/rv32i_test")
    ) u3 (
        .clk            (clk), 
        .funct3         (funct3), 
        .dmem_wren      (dmem_wren), 
        .dmem_address   (dmem_address), 
        .dmem_data_in   (dmem_data_in), 
        .imem_address   (imem_address), 
        .imem_data_out  (imem_data_out), 
        .dmem_data_out  (dmem_data_out), 
        .reset          (reset), 
        .led            (led), 
        .red            (red), 
        .green          (green), 
        .blue           (blue)
    );

    assign LED = ~led;
    assign RGB_R = ~red;
    assign RGB_G = ~green;
    assign RGB_B = ~blue;

endmodule