/*
 *  Program Counter
 *  
 *  Program Counter for RISC-V Processor
 */